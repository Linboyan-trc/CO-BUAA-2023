module IM(
    input [31:0] PC,
    output [31:0] Ins
);
    //ROM
    reg [31:0] IMdeROM [0:4095];

    // //载入指令
    // initial begin
    //     $readmemh("code.txt",IMdeROM);
    // end
    //vscode专用载入指令
    initial begin
        IMdeROM[0]<=32'h34010006;
        IMdeROM[1]<=32'h34020003;
        IMdeROM[2]<=32'h34030005;
        IMdeROM[3]<=32'h34040009;
        IMdeROM[4]<=32'h3405000c;
        IMdeROM[5]<=32'h34060005;
        IMdeROM[6]<=32'h34070009;
        IMdeROM[7]<=32'h3408000a;
        IMdeROM[8]<=32'h34090005;
        IMdeROM[9]<=32'h340a0004;
        IMdeROM[10]<=32'h340b0004;
        IMdeROM[11]<=32'h340c0004;
        IMdeROM[12]<=32'h340d000a;
        IMdeROM[13]<=32'h340e0004;
        IMdeROM[14]<=32'h340f0006;
        IMdeROM[15]<=32'h34100005;
        IMdeROM[16]<=32'h34110007;
        IMdeROM[17]<=32'h3412000b;
        IMdeROM[18]<=32'h34130006;
        IMdeROM[19]<=32'h3414000c;
        IMdeROM[20]<=32'h34150003;
        IMdeROM[21]<=32'h34160003;
        IMdeROM[22]<=32'h34170004;
        IMdeROM[23]<=32'h3418000a;
        IMdeROM[24]<=32'h34190008;
        IMdeROM[25]<=32'h341a000a;
        IMdeROM[26]<=32'h341b0005;
        IMdeROM[27]<=32'h341c0006;
        IMdeROM[28]<=32'h341d0004;
        IMdeROM[29]<=32'h341e000a;
        IMdeROM[30]<=32'h347900ed;
        IMdeROM[31]<=32'h0c000c24;
        IMdeROM[32]<=32'h00000000;
        IMdeROM[33]<=32'h3479017b;
        IMdeROM[34]<=32'h0c000c4c;
        IMdeROM[35]<=32'h00000000;
        IMdeROM[36]<=32'h3c0601be;
        IMdeROM[37]<=32'h340b0008;
        IMdeROM[38]<=32'h8d630024;
        IMdeROM[39]<=32'h0004e020;
        IMdeROM[40]<=32'h368e012c;
        IMdeROM[41]<=32'h341d0010;
        IMdeROM[42]<=32'h8fb90098;
        IMdeROM[43]<=32'h3c1d0067;
        IMdeROM[44]<=32'h00000000;
        IMdeROM[45]<=32'h02924020;
        IMdeROM[46]<=32'h3c1e0055;
        IMdeROM[47]<=32'h03aef022;
        IMdeROM[48]<=32'h34150095;
        IMdeROM[49]<=32'h359f01c4;
        IMdeROM[50]<=32'h34170004;
        IMdeROM[51]<=32'haeeb0020;
        IMdeROM[52]<=32'h00000000;
        IMdeROM[53]<=32'h00000000;
        IMdeROM[54]<=32'h3c040008;
        IMdeROM[55]<=32'h341e000c;
        IMdeROM[56]<=32'hafcc0028;
        IMdeROM[57]<=32'h34010010;
        IMdeROM[58]<=32'h8c370040;
        IMdeROM[59]<=32'h347c0164;
        IMdeROM[60]<=32'h34070010;
        IMdeROM[61]<=32'h8ce8008c;
        IMdeROM[62]<=32'h3c010023;
        IMdeROM[63]<=32'h341c0010;
        IMdeROM[64]<=32'h8f870084;
        IMdeROM[65]<=32'h363b00b6;
        IMdeROM[66]<=32'h016d4020;
        IMdeROM[67]<=32'h343c00e4;
        IMdeROM[68]<=32'h36bf00d8;
        IMdeROM[69]<=32'h3c1a009c;
        IMdeROM[70]<=32'h01473822;
        IMdeROM[71]<=32'h34160014;
        IMdeROM[72]<=32'haece008c;
        IMdeROM[73]<=32'h3c020101;
        IMdeROM[74]<=32'h1361ffd6;
        IMdeROM[75]<=32'h00000000;
        IMdeROM[76]<=32'h0c000c51;
        IMdeROM[77]<=32'h00000000;
        IMdeROM[78]<=32'h3c1b00af;
        IMdeROM[79]<=32'h0c000c7c;
        IMdeROM[80]<=32'h00000000;
        IMdeROM[81]<=32'h35d1001f;
        IMdeROM[82]<=32'h00000000;
        IMdeROM[83]<=32'h340d0014;
        IMdeROM[84]<=32'hadb00010;
        IMdeROM[85]<=32'h3411000c;
        IMdeROM[86]<=32'h8e2d0038;
        IMdeROM[87]<=32'h361d0156;
        IMdeROM[88]<=32'h340e0014;
        IMdeROM[89]<=32'h8dd70078;
        IMdeROM[90]<=32'h00000000;
        IMdeROM[91]<=32'h00000000;
        IMdeROM[92]<=32'h004a7820;
        IMdeROM[93]<=32'h37e8003a;
        IMdeROM[94]<=32'h009ce022;
        IMdeROM[95]<=32'h3c1b018e;
        IMdeROM[96]<=32'h039ab822;
        IMdeROM[97]<=32'h34010018;
        IMdeROM[98]<=32'hac3d0060;
        IMdeROM[99]<=32'h3c1b0037;
        IMdeROM[100]<=32'h34100008;
        IMdeROM[101]<=32'h8e040028;
        IMdeROM[102]<=32'h34100014;
        IMdeROM[103]<=32'h8e0d000c;
        IMdeROM[104]<=32'h012bb820;
        IMdeROM[105]<=32'h34110008;
        IMdeROM[106]<=32'h8e270084;
        IMdeROM[107]<=32'h340a000c;
        IMdeROM[108]<=32'had57005c;
        IMdeROM[109]<=32'h00000000;
        IMdeROM[110]<=32'h01952022;
        IMdeROM[111]<=32'h02999020;
        IMdeROM[112]<=32'h34100018;
        IMdeROM[113]<=32'h8e110014;
        IMdeROM[114]<=32'h00000000;
        IMdeROM[115]<=32'h341e0004;
        IMdeROM[116]<=32'hafcf0078;
        IMdeROM[117]<=32'h34e30191;
        IMdeROM[118]<=32'h00892020;
        IMdeROM[119]<=32'h34060010;
        IMdeROM[120]<=32'h8cd70000;
        IMdeROM[121]<=32'h00000000;
        IMdeROM[122]<=32'h1026ffd3;
        IMdeROM[123]<=32'h00000000;
        IMdeROM[124]<=32'h0c000c81;
        IMdeROM[125]<=32'h00000000;
        IMdeROM[126]<=32'h00000000;
        IMdeROM[127]<=32'h0c000ca5;
        IMdeROM[128]<=32'h00000000;
        IMdeROM[129]<=32'h375400b1;
        IMdeROM[130]<=32'h021be022;
        IMdeROM[131]<=32'h01881020;
        IMdeROM[132]<=32'h34080014;
        IMdeROM[133]<=32'h8d1b002c;
        IMdeROM[134]<=32'h349f011c;
        IMdeROM[135]<=32'h022a8822;
        IMdeROM[136]<=32'h0372b022;
        IMdeROM[137]<=32'h34080014;
        IMdeROM[138]<=32'h8d1b0040;
        IMdeROM[139]<=32'h340c014a;
        IMdeROM[140]<=32'h341c0014;
        IMdeROM[141]<=32'haf9900a0;
        IMdeROM[142]<=32'h00000000;
        IMdeROM[143]<=32'h37df019d;
        IMdeROM[144]<=32'h3c040128;
        IMdeROM[145]<=32'h3c0400a3;
        IMdeROM[146]<=32'h3c010196;
        IMdeROM[147]<=32'h00000000;
        IMdeROM[148]<=32'h3c1001c0;
        IMdeROM[149]<=32'h01c38822;
        IMdeROM[150]<=32'h00d1d020;
        IMdeROM[151]<=32'h0057d822;
        IMdeROM[152]<=32'h034f3022;
        IMdeROM[153]<=32'h3c060097;
        IMdeROM[154]<=32'h34020014;
        IMdeROM[155]<=32'hac480034;
        IMdeROM[156]<=32'h0276f022;
        IMdeROM[157]<=32'h3c170138;
        IMdeROM[158]<=32'h34160004;
        IMdeROM[159]<=32'h8ec50094;
        IMdeROM[160]<=32'h00000000;
        IMdeROM[161]<=32'h34d40080;
        IMdeROM[162]<=32'h3c0b0162;
        IMdeROM[163]<=32'h1257ffda;
        IMdeROM[164]<=32'h00000000;
        IMdeROM[165]<=32'h13ee0028;
        IMdeROM[166]<=32'h00000000;
        IMdeROM[167]<=32'h00000000;
        IMdeROM[168]<=32'h37fd0028;
        IMdeROM[169]<=32'h017ea020;
        IMdeROM[170]<=32'h0023d820;
        IMdeROM[171]<=32'h350e0012;
        IMdeROM[172]<=32'h3419000c;
        IMdeROM[173]<=32'haf23001c;
        IMdeROM[174]<=32'h01687820;
        IMdeROM[175]<=32'h341a0010;
        IMdeROM[176]<=32'h8f450064;
        IMdeROM[177]<=32'h34180008;
        IMdeROM[178]<=32'haf0a0044;
        IMdeROM[179]<=32'h0363e822;
        IMdeROM[180]<=32'h027d8022;
        IMdeROM[181]<=32'h00fc4820;
        IMdeROM[182]<=32'h34010014;
        IMdeROM[183]<=32'hac380094;
        IMdeROM[184]<=32'h00000000;
        IMdeROM[185]<=32'h02ade020;
        IMdeROM[186]<=32'h3c0700a2;
        IMdeROM[187]<=32'h3c0501b9;
        IMdeROM[188]<=32'h3c1a0160;
        IMdeROM[189]<=32'h00000000;
        IMdeROM[190]<=32'h007d1020;
        IMdeROM[191]<=32'h3c18018d;
        IMdeROM[192]<=32'h353801c2;
        IMdeROM[193]<=32'h006dd020;
        IMdeROM[194]<=32'h341e000c;
        IMdeROM[195]<=32'hafca008c;
        IMdeROM[196]<=32'h34050014;
        IMdeROM[197]<=32'hacb00014;
        IMdeROM[198]<=32'h3413000c;
        IMdeROM[199]<=32'hae6b0004;
        IMdeROM[200]<=32'h00000000;
        IMdeROM[201]<=32'h032d5820;
        IMdeROM[202]<=32'h34190014;
        IMdeROM[203]<=32'haf3c0020;
        IMdeROM[204]<=32'h10480001;
        IMdeROM[205]<=32'h00000000;
        IMdeROM[206]<=32'h36dc01a8;
        IMdeROM[207]<=32'h341d000c;
        IMdeROM[208]<=32'h8faa002c;
        IMdeROM[209]<=32'h00764020;
        IMdeROM[210]<=32'h34130010;
        IMdeROM[211]<=32'hae680060;
        IMdeROM[212]<=32'h36c20015;
        IMdeROM[213]<=32'h0244c822;
        IMdeROM[214]<=32'h34010014;
        IMdeROM[215]<=32'h8c250010;
        IMdeROM[216]<=32'h352701bb;
        IMdeROM[217]<=32'h03196820;
        IMdeROM[218]<=32'h34180008;
        IMdeROM[219]<=32'haf000004;
        IMdeROM[220]<=32'h3c1b0186;
        IMdeROM[221]<=32'h34130004;
        IMdeROM[222]<=32'h8e6600a0;
        IMdeROM[223]<=32'h00946020;
        IMdeROM[224]<=32'h03bd3820;
        IMdeROM[225]<=32'h00000000;
        IMdeROM[226]<=32'hac180054;
        IMdeROM[227]<=32'h37a1001c;
        IMdeROM[228]<=32'h00000000;
        IMdeROM[229]<=32'h34090010;
        IMdeROM[230]<=32'had250034;
        IMdeROM[231]<=32'h0082b822;
        IMdeROM[232]<=32'h0249b822;
        IMdeROM[233]<=32'h350900bb;
        IMdeROM[234]<=32'h03a5c020;
        IMdeROM[235]<=32'h3c14002f;
        IMdeROM[236]<=32'h37730057;
        IMdeROM[237]<=32'h3c05017d;
        IMdeROM[238]<=32'h00cfb822;
        IMdeROM[239]<=32'h353300f8;
        IMdeROM[240]<=32'h027ac022;
        IMdeROM[241]<=32'h11e30001;
        IMdeROM[242]<=32'h00000000;
        IMdeROM[243]<=32'h340f000c;
        IMdeROM[244]<=32'h8df50074;
        IMdeROM[245]<=32'h017cd820;
        IMdeROM[246]<=32'h340b0004;
        IMdeROM[247]<=32'had6e0078;
        IMdeROM[248]<=32'h00aac022;
        IMdeROM[249]<=32'h341a0010;
        IMdeROM[250]<=32'h8f590080;
        IMdeROM[251]<=32'h00000000;
        IMdeROM[252]<=32'h00000000;
        IMdeROM[253]<=32'h00000000;
        IMdeROM[254]<=32'h00000000;
        IMdeROM[255]<=32'h01359820;
        IMdeROM[256]<=32'h34480010;
        IMdeROM[257]<=32'h00000000;
        IMdeROM[258]<=32'h3415000c;
        IMdeROM[259]<=32'h8ea10000;
        IMdeROM[260]<=32'h00000000;
        IMdeROM[261]<=32'h00f01022;
        IMdeROM[262]<=32'h01ff2022;
        IMdeROM[263]<=32'h34130004;
        IMdeROM[264]<=32'h8e760010;
        IMdeROM[265]<=32'h3c1a0127;
        IMdeROM[266]<=32'h3c150171;
        IMdeROM[267]<=32'h0265c822;
        IMdeROM[268]<=32'h02c17020;
        IMdeROM[269]<=32'h34010008;
        IMdeROM[270]<=32'h8c2f0084;
        IMdeROM[271]<=32'h341e0008;
        IMdeROM[272]<=32'h8fc30018;
        IMdeROM[273]<=32'h3401000c;
        IMdeROM[274]<=32'hac2d00a0;
        IMdeROM[275]<=32'h34160010;
        IMdeROM[276]<=32'h8ec6009c;
        IMdeROM[277]<=32'h34190004;
        IMdeROM[278]<=32'h8f3e0084;
        IMdeROM[279]<=32'h34150014;
        IMdeROM[280]<=32'haeb50064;
        IMdeROM[281]<=32'h34140008;
        IMdeROM[282]<=32'hae98007c;
        IMdeROM[283]<=32'h340d0004;
        IMdeROM[284]<=32'hadb90084;
        IMdeROM[285]<=32'h122c0001;
        IMdeROM[286]<=32'h00000000;
        IMdeROM[287]<=32'h3c0e00e4;
        IMdeROM[288]<=32'h34c60117;
        IMdeROM[289]<=32'h00000000;
        IMdeROM[290]<=32'h022d5822;
        IMdeROM[291]<=32'h360700cd;
        IMdeROM[292]<=32'h00000000;
        IMdeROM[293]<=32'h039b2022;
        IMdeROM[294]<=32'h340a0014;
        IMdeROM[295]<=32'h8d45004c;
        IMdeROM[296]<=32'h3c1c0016;
        IMdeROM[297]<=32'h340f0018;
        IMdeROM[298]<=32'h8def0090;
        IMdeROM[299]<=32'h34050014;
        IMdeROM[300]<=32'h8cac0038;
        IMdeROM[301]<=32'hac130074;
        IMdeROM[302]<=32'h002a4020;
        IMdeROM[303]<=32'h35690028;
        IMdeROM[304]<=32'h3c07019b;
        IMdeROM[305]<=32'h3c1200e0;
        IMdeROM[306]<=32'h36d70181;
        IMdeROM[307]<=32'h34110008;
        IMdeROM[308]<=32'hae3e008c;
        IMdeROM[309]<=32'h34150010;
        IMdeROM[310]<=32'haebe0050;
    end

    //输出Ins
    wire [31:0]tempPC;
    assign tempPC=PC-32'h0000_3000;
    assign Ins=IMdeROM[tempPC[13:2]];
endmodule