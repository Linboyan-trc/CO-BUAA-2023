module testclk(input a);
    
endmodule